`include "cu.sv"
`include "decode.sv"
`include "exec.sv"
`include "fetch.sv"
`include "mem.sv"
`include "pc.sv"
`include "pipeline_dec.sv"
`include "pipeline_ex.sv"
`include "pipeline_fetch.sv"
`include "pipeline_mem.sv"
`include "regfile.sv"










