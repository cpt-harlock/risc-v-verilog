`define FETCH_SEL_PC 2'b00
`define FETCH_SEL_BRANCH 2'b01
`define FETCH_SEL_NOP 2'b10
`define FETCH_SEL_NOP 2'b10
`define NOP_INSTRUCTION 32'b0000000_00000_00000_000_00000_0110011
`define NOP_INSTRUCTION_OPCODE 32'b0110011
`define NOP_INSTRUCTION_RD 5'b00000
`define NOP_INSTRUCTION_FUNCT3 3'b000
`define NOP_INSTRUCTION_FUNCT7 7'b0000000
`define NOP_INSTRUCTION_RS1 5'b00000
`define NOP_INSTRUCTION_RS1_DATA 32'b00000
`define NOP_INSTRUCTION_RS2 5'b00000
`define NOP_INSTRUCTION_RS2_DATA 32'b00000
`define NOP_INSTRUCTION_IMM 32'b0
`define NOP_INSTRUCTION_PC 32'b0
`define DATA_MEM_SIZE 2**10
`define INSTRUCTIONS_MEM_SIZE 2**8

`define R 3'b000
`define I 3'b001
`define S 3'b010
`define B 3'b011 
`define U 3'b100
`define J 3'b101
`define WRONG_INSTRUCTION_TYPE 3'b111