`define LB 'b0000011_000_x
`define LH 'b0000011_001_x
`define LW 'b0000011_010_x
`define LBU 'b0000011_100_x
`define LHU 'b0000011_101_x
`define ADDI 'b0010011_000_x
`define SLLI 'b0010011_001_0
`define SLTI 'b0010011_010_x
`define SLTIU 'b0010011_011_x
`define XORI 'b0010011_100_x
`define SRLI 'b0010011_101_0
`define SRAI 'b0010011_101_1
`define ORI 'b0010011_110_1
`define ANDI 'b0010011_111_1
`define AUIPC 'b0010111_xxx_x
`define SB 'b0100011_000_x
`define SH 'b0100011_001_x
`define SW 'b0100011_010_x
`define ADD 'b0110011_000_0
`define SUB 'b0110011_000_1
`define SLL 'b0110011_001_0
`define SLT 'b0110011_010_0
`define SLTU 'b0110011_011_0
`define XOR 'b0110011_100_0
`define SRL 'b0110011_101_0
`define SRA 'b0110011_101_1
`define OR 'b0110011_110_0
`define AND 'b0110011_111_0
`define LUI 'b0110111_xxx_x
`define BEQ 'b1100011_000_x
`define BNE 'b1100011_001_x
`define BLT 'b1100011_100_x
`define BGE 'b1100011_101_x
`define BLTU 'b1100011_110_x
`define BGEU 'b1100011_111_x
`define JALR 'b1100111_000_x
`define JAL 'b1101111_xxx_x

