`define LB 'b0000011_000_? //OK
`define LH 'b0000011_001_? //OK 
`define LW 'b0000011_010_? //OK 
`define LBU 'b0000011_100_? // OK 
`define LHU 'b0000011_101_? // OK 
`define ADDI 'b0010011_000_? // OK
`define SLLI 'b0010011_001_0 // OK 
`define SLTI 'b0010011_010_? // OK 
`define SLTIU 'b0010011_011_? // OK 
`define XORI 'b0010011_100_? // OK 
`define SRLI 'b0010011_101_0 // OK 
`define SRAI 'b0010011_101_1 // OK 
`define ORI 'b0010011_110_? // OK 
`define ANDI 'b0010011_111_? // OK 
`define AUIPC 'b0010111_???_? // OK 
`define SB 'b0100011_000_? // OK 
`define SH 'b0100011_001_? // OK 
`define SW 'b0100011_010_? // OK 
`define ADD 'b0110011_000_0 //OK
`define SUB 'b0110011_000_1 //OK
`define SLL 'b0110011_001_0 // OK 
`define SLT 'b0110011_010_0 // OK 
`define SLTU 'b0110011_011_0 // OK 
`define XOR 'b0110011_100_0 // OK 
`define SRL 'b0110011_101_0 // OK 
`define SRA 'b0110011_101_1 // OK 
`define OR 'b0110011_110_0 // OK 
`define AND 'b0110011_111_0 // OK
`define LUI 'b0110111_???_? // OK 
`define BEQ 'b1100011_000_? // OK 
`define BNE 'b1100011_001_? // OK 
`define BLT 'b1100011_100_? // OK 
`define BGE 'b1100011_101_? // OK 
`define BLTU 'b1100011_110_? // OK 
`define BGEU 'b1100011_111_? // OK 
`define JALR 'b1100111_000_? // OK 
`define JAL 'b1101111_???_? // OK 

