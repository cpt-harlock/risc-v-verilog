`define LB 'b0000011_000_?
`define LH 'b0000011_001_?
`define LW 'b0000011_010_?
`define LBU 'b0000011_100_?
`define LHU 'b0000011_101_?
`define ADDI 'b0010011_000_?
`define SLLI 'b0010011_001_0
`define SLTI 'b0010011_010_?
`define SLTIU 'b0010011_011_?
`define XORI 'b0010011_100_?
`define SRLI 'b0010011_101_0
`define SRAI 'b0010011_101_1
`define ORI 'b0010011_110_1
`define ANDI 'b0010011_111_1
`define AUIPC 'b0010111_???_?
`define SB 'b0100011_000_?
`define SH 'b0100011_001_?
`define SW 'b0100011_010_?
`define ADD 'b0110011_000_0
`define SUB 'b0110011_000_1
`define SLL 'b0110011_001_0
`define SLT 'b0110011_010_0
`define SLTU 'b0110011_011_0
`define XOR 'b0110011_100_0
`define SRL 'b0110011_101_0
`define SRA 'b0110011_101_1
`define OR 'b0110011_110_0
`define AND 'b0110011_111_0
`define LUI 'b0110111_???_?
`define BEQ 'b1100011_000_?
`define BNE 'b1100011_001_?
`define BLT 'b1100011_100_?
`define BGE 'b1100011_101_?
`define BLTU 'b1100011_110_?
`define BGEU 'b1100011_111_?
`define JALR 'b1100111_000_?
`define JAL 'b1101111_???_?

